--
-- VHDL Architecture PTR3_HVPS_lib.HVPS_I2C.beh
--
-- Created:
--          by - nort.UNKNOWN (NORT-XPS14)
--          at - 11:08:55 11/ 8/2016
--
-- using Mentor Graphics HDL Designer(TM) 2013.1b (Build 2)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY aio_i2c IS
   PORT( 
      rst       : IN     std_ulogic;
      wb_adr_i  : IN     std_logic_vector (2 DOWNTO 0);
      wb_cyc_i  : IN     std_logic;
      wb_dat_i  : IN     std_logic_vector (7 DOWNTO 0);
      wb_stb_i  : IN     std_logic;
      wb_we_i   : IN     std_logic;
      scl_pad_i    : IN  std_logic;
      scl_pad_o    : OUT std_logic;
      scl_padoen_o : OUT std_logic;
      sda_pad_i    : IN  std_logic;
      sda_pad_o    : OUT std_logic;
      sda_padoen_o : OUT std_logic;
      wb_ack_o  : OUT    std_logic;
      wb_dat_o  : OUT    std_logic_vector (7 DOWNTO 0);
      wb_inta_o : OUT    std_logic;
      clk       : IN     std_ulogic
   );

-- Declarations

END aio_i2c ;

--
ARCHITECTURE beh OF aio_i2c IS

   COMPONENT i2c_master_top
      GENERIC (
         ARST_LVL : std_logic := '0'
      );
      PORT (
         wb_clk_i     : IN     std_logic;
         wb_rst_i     : IN     std_logic;
         arst_i       : IN     std_logic;
         wb_adr_i     : IN     std_logic_vector(2 downto 0);
         wb_dat_i     : IN     std_logic_vector(7 downto 0);
         wb_dat_o     : OUT    std_logic_vector(7 downto 0);
         wb_we_i      : IN     std_logic;
         wb_stb_i     : IN     std_logic;
         wb_cyc_i     : IN     std_logic;
         wb_ack_o     : OUT    std_logic;
         wb_inta_o    : OUT    std_logic;
         scl_pad_i    : IN     std_logic;
         scl_pad_o    : OUT    std_logic;
         scl_padoen_o : OUT    std_logic;
         sda_pad_i    : IN     std_logic;
         sda_pad_o    : OUT    std_logic;
         sda_padoen_o : OUT    std_logic
      );
   END COMPONENT;
BEGIN
   --  hds hds_inst
   i2c_master : i2c_master_top
      GENERIC MAP (
         ARST_LVL => '0'
      )
      PORT MAP (
         wb_clk_i     => clk,
         wb_rst_i     => rst,
         arst_i       => '1',
         wb_adr_i     => wb_adr_i,
         wb_dat_i     => wb_dat_i,
         wb_dat_o     => wb_dat_o,
         wb_we_i      => wb_we_i,
         wb_stb_i     => wb_stb_i,
         wb_cyc_i     => wb_cyc_i,
         wb_ack_o     => wb_ack_o,
         wb_inta_o    => wb_inta_o,
         scl_pad_i    => scl_pad_i,
         scl_pad_o    => scl_pad_o,
         scl_padoen_o => scl_padoen_o,
         sda_pad_i    => sda_pad_i,
         sda_pad_o    => sda_pad_o,
         sda_padoen_o => sda_padoen_o
      );
END ARCHITECTURE beh;

